avg-delay,mode,benchmark,iteration,tail-latency
0.1,cpu,imc,1,3871.184502
0.1,cpu,dig,1,624.000294
0.1,cpu,face,1,0
0.1,cpu,ner,1,183.806748
0.1,shared_gpu,imc,1,33.725339
0.1,shared_gpu,dig,1,6.091226
0.1,shared_gpu,face,1,233.065173
0.1,shared_gpu,ner,1,48.191989
0.1,dedicated_gpu,imc,1,108.429013
0.1,dedicated_gpu,dig,1,11.953061
0.1,dedicated_gpu,face,1,189.762973
0.1,dedicated_gpu,ner,1,75.010397
0.25,cpu,imc,1,1627.965924
0.25,cpu,dig,1,159.954881
0.25,cpu,face,1,5165.36153
0.25,cpu,ner,1,67.590353
0.25,shared_gpu,imc,1,23.761833
0.25,shared_gpu,dig,1,2.887623
0.25,shared_gpu,face,1,103.452175
0.25,shared_gpu,ner,1,55.648816
0.25,dedicated_gpu,imc,1,21.273042
0.25,dedicated_gpu,dig,1,8.271139
0.25,dedicated_gpu,face,1,99.893979
0.25,dedicated_gpu,ner,1,5.02901
0.5,cpu,imc,1,1956.477337
0.5,cpu,dig,1,198.917049
0.5,cpu,face,1,5459.928996
0.5,cpu,ner,1,178.405543
0.5,shared_gpu,imc,1,26.961382
0.5,shared_gpu,dig,1,11.178933
0.5,shared_gpu,face,1,91.006985
0.5,shared_gpu,ner,1,42.114491
0.5,dedicated_gpu,imc,1,13.68898
0.5,dedicated_gpu,dig,1,12.687876
0.5,dedicated_gpu,face,1,93.134251
0.5,dedicated_gpu,ner,1,12.965899
1,cpu,imc,1,843.893261
1,cpu,dig,1,125.779544
1,cpu,face,1,2018.638855
1,cpu,ner,1,54.656847
1,shared_gpu,imc,1,18.803183
1,shared_gpu,dig,1,6.948829
1,shared_gpu,face,1,35.652463
1,shared_gpu,ner,1,20.949192
1,dedicated_gpu,imc,1,13.649125
1,dedicated_gpu,dig,1,5.875575
1,dedicated_gpu,face,1,37.083593
1,dedicated_gpu,ner,1,21.443668
0.25,cpu,imc,2,1511.605824
0.25,cpu,dig,2,113.210744
0.25,cpu,face,2,5287.946859
0.25,cpu,ner,2,64.430665
0.25,shared_gpu,imc,2,19.904847
0.25,shared_gpu,dig,2,4.927728
0.25,shared_gpu,face,2,100.207283
0.25,shared_gpu,ner,2,75.576379
0.25,dedicated_gpu,imc,2,29.889955
0.25,dedicated_gpu,dig,2,10.582027
0.25,dedicated_gpu,face,2,110.084609
0.25,dedicated_gpu,ner,2,31.619233
1,cpu,imc,2,1009.469916
1,cpu,dig,2,74.676303
1,cpu,face,2,2179.385198
1,cpu,ner,2,75.539247
1,shared_gpu,imc,2,10.143573
1,shared_gpu,dig,2,4.185463
1,shared_gpu,face,2,34.245976
1,shared_gpu,ner,2,25.354584
1,dedicated_gpu,imc,2,12.344335
1,dedicated_gpu,dig,2,5.274144
1,dedicated_gpu,face,2,32.094453
1,dedicated_gpu,ner,2,9.638261
0.5,cpu,imc,2,2277.753796
0.5,cpu,dig,2,158.703544
0.5,cpu,face,2,5472.705603
0.5,cpu,ner,2,93.616017
0.5,shared_gpu,imc,2,29.97071
0.5,shared_gpu,dig,2,4.20552
0.5,shared_gpu,face,2,101.82666
0.5,shared_gpu,ner,2,45.480191
0.5,dedicated_gpu,imc,2,0
0.5,dedicated_gpu,dig,2,4.078233
0.5,dedicated_gpu,face,2,0
0.5,dedicated_gpu,ner,2,0
0.1,cpu,imc,2,3479.524377
0.1,cpu,dig,2,246.808776
0.1,cpu,face,2,0
0.1,cpu,ner,2,99.775846
0.1,shared_gpu,imc,2,32.419586
0.1,shared_gpu,dig,2,5.302847
0.1,shared_gpu,face,2,191.832184
0.1,shared_gpu,ner,2,54.879148
0.1,dedicated_gpu,imc,2,30.13082
0.1,dedicated_gpu,dig,2,6.913026
0.1,dedicated_gpu,face,2,207.147694
0.1,dedicated_gpu,ner,2,128.605272
0.25,cpu,imc,3,1538.65726
0.25,cpu,dig,3,244.154393
0.25,cpu,face,3,5263.4584
0.25,cpu,ner,3,104.084386
0.25,shared_gpu,imc,3,23.411838
0.25,shared_gpu,dig,3,11.569307
0.25,shared_gpu,face,3,99.862579
0.25,shared_gpu,ner,3,77.939351
0.25,dedicated_gpu,imc,3,25.681636
0.25,dedicated_gpu,dig,3,8.409553
0.25,dedicated_gpu,face,3,106.410647
0.25,dedicated_gpu,ner,3,53.548586
0.1,cpu,imc,3,3658.696133
0.1,cpu,dig,3,288.671659
0.1,cpu,face,3,0
0.1,cpu,ner,3,119.873497
0.1,shared_gpu,imc,3,47.46605
0.1,shared_gpu,dig,3,6.544742
0.1,shared_gpu,face,3,191.785026
0.1,shared_gpu,ner,3,187.524075
0.1,dedicated_gpu,imc,3,110.675786
0.1,dedicated_gpu,dig,3,6.835985
0.1,dedicated_gpu,face,3,198.199583
0.1,dedicated_gpu,ner,3,99.561388
0.5,cpu,imc,3,1793.629246
0.5,cpu,dig,3,122.566039
0.5,cpu,face,3,5637.964938
0.5,cpu,ner,3,87.967082
0.5,shared_gpu,imc,3,25.046936
0.5,shared_gpu,dig,3,14.36606
0.5,shared_gpu,face,3,96.320423
0.5,shared_gpu,ner,3,9.868032
0.5,dedicated_gpu,imc,3,20.110421
0.5,dedicated_gpu,dig,3,9.555388
0.5,dedicated_gpu,face,3,71.983793
0.5,dedicated_gpu,ner,3,8.558422
1,cpu,imc,3,888.764783
1,cpu,dig,3,78.479271
1,cpu,face,3,1946.109111
1,cpu,ner,3,130.783615
1,shared_gpu,imc,3,18.410696
1,shared_gpu,dig,3,10.453254
1,shared_gpu,face,3,33.792239
1,shared_gpu,ner,3,4.559507
1,dedicated_gpu,imc,3,0
1,dedicated_gpu,dig,3,2.926855
1,dedicated_gpu,face,3,0
1,dedicated_gpu,ner,3,0
1,cpu,imc,4,918.29335
1,cpu,dig,4,145.2275
1,cpu,face,4,2119.004038
1,cpu,ner,4,75.955551
1,shared_gpu,imc,4,10.144468
1,shared_gpu,dig,4,7.65175
1,shared_gpu,face,4,34.535427
1,shared_gpu,ner,4,19.472103
1,dedicated_gpu,imc,4,13.372569
1,dedicated_gpu,dig,4,4.02845
1,dedicated_gpu,face,4,37.599178
1,dedicated_gpu,ner,4,19.561033
0.25,cpu,imc,4,2089.669836
0.25,cpu,dig,4,200.444424
0.25,cpu,face,4,6175.207406
0.25,cpu,ner,4,79.340327
0.25,shared_gpu,imc,4,18.984738
0.25,shared_gpu,dig,4,6.071759
0.25,shared_gpu,face,4,108.509043
0.25,shared_gpu,ner,4,61.406739
0.25,dedicated_gpu,imc,4,27.426634
0.25,dedicated_gpu,dig,4,5.858788
0.25,dedicated_gpu,face,4,99.898957
0.25,dedicated_gpu,ner,4,12.15678
0.5,cpu,imc,4,1646.357102
0.5,cpu,dig,4,459.096676
0.5,cpu,face,4,5337.234095
0.5,cpu,ner,4,75.241502
0.5,shared_gpu,imc,4,15.412495
0.5,shared_gpu,dig,4,11.122773
0.5,shared_gpu,face,4,93.688885
0.5,shared_gpu,ner,4,52.222145
0.5,dedicated_gpu,imc,4,23.42565
0.5,dedicated_gpu,dig,4,7.722443
0.5,dedicated_gpu,face,4,96.335959
0.5,dedicated_gpu,ner,4,13.09507
0.1,cpu,imc,4,3481.362364
0.1,cpu,dig,4,347.53239
0.1,cpu,face,4,0
0.1,cpu,ner,4,59.679606
0.1,shared_gpu,imc,4,46.203756
0.1,shared_gpu,dig,4,16.914212
0.1,shared_gpu,face,4,196.299042
0.1,shared_gpu,ner,4,63.933737
0.1,dedicated_gpu,imc,4,40.883164
0.1,dedicated_gpu,dig,4,4.774283
0.1,dedicated_gpu,face,4,132.1263
0.1,dedicated_gpu,ner,4,8.022389
1,cpu,imc,5,660.189817
1,cpu,dig,5,112.433975
1,cpu,face,5,1812.865637
1,cpu,ner,5,47.195675
1,shared_gpu,imc,5,9.229565
1,shared_gpu,dig,5,3.524854
1,shared_gpu,face,5,35.098196
1,shared_gpu,ner,5,23.480272
1,dedicated_gpu,imc,5,14.077799
1,dedicated_gpu,dig,5,5.488028
1,dedicated_gpu,face,5,37.958923
1,dedicated_gpu,ner,5,23.449748
0.25,cpu,imc,5,1644.301092
0.25,cpu,dig,5,254.529966
0.25,cpu,face,5,5145.587763
0.25,cpu,ner,5,52.479582
0.25,shared_gpu,imc,5,20.011329
0.25,shared_gpu,dig,5,15.464541
0.25,shared_gpu,face,5,121.496455
0.25,shared_gpu,ner,5,72.968875
0.25,dedicated_gpu,imc,5,26.7879
0.25,dedicated_gpu,dig,5,7.800166
0.25,dedicated_gpu,face,5,107.415009
0.25,dedicated_gpu,ner,5,41.23415
0.5,cpu,imc,5,2055.031274
0.5,cpu,dig,5,230.457288
0.5,cpu,face,5,5728.896797
0.5,cpu,ner,5,117.319363
0.5,shared_gpu,imc,5,17.976476
0.5,shared_gpu,dig,5,6.566833
0.5,shared_gpu,face,5,93.275509
0.5,shared_gpu,ner,5,55.679354
0.5,dedicated_gpu,imc,5,17.505946
0.5,dedicated_gpu,dig,5,6.311598
0.5,dedicated_gpu,face,5,95.04387
0.5,dedicated_gpu,ner,5,43.389153
0.1,cpu,imc,5,3370.579561
0.1,cpu,dig,5,372.197043
0.1,cpu,face,5,0
0.1,cpu,ner,5,104.127821
0.1,shared_gpu,imc,5,38.040309
0.1,shared_gpu,dig,5,26.45805
0.1,shared_gpu,face,5,184.983995
0.1,shared_gpu,ner,5,175.963032
0.1,dedicated_gpu,imc,5,43.081167
0.1,dedicated_gpu,dig,5,11.758003
0.1,dedicated_gpu,face,5,194.773421
0.1,dedicated_gpu,ner,5,50.68696
1,cpu,imc,6,802.37376
1,cpu,dig,6,210.705701
1,cpu,face,6,2102.655107
1,cpu,ner,6,87.32119
1,shared_gpu,imc,6,12.297483
1,shared_gpu,dig,6,6.507823
1,shared_gpu,face,6,33.786755
1,shared_gpu,ner,6,12.07908
1,dedicated_gpu,imc,6,12.504939
1,dedicated_gpu,dig,6,6.329774
1,dedicated_gpu,face,6,36.886836
1,dedicated_gpu,ner,6,18.29168
0.25,cpu,imc,6,1717.804913
0.25,cpu,dig,6,162.624782
0.25,cpu,face,6,5261.402429
0.25,cpu,ner,6,42.447818
0.25,shared_gpu,imc,6,18.678914
0.25,shared_gpu,dig,6,4.70887
0.25,shared_gpu,face,6,101.744966
0.25,shared_gpu,ner,6,62.424631
0.25,dedicated_gpu,imc,6,24.078957
0.25,dedicated_gpu,dig,6,5.642869
0.25,dedicated_gpu,face,6,101.960212
0.25,dedicated_gpu,ner,6,32.629106
0.1,cpu,imc,6,3471.036626
0.1,cpu,dig,6,228.590725
0.1,cpu,face,6,0
0.1,cpu,ner,6,80.524516
0.1,shared_gpu,imc,6,158.909514
0.1,shared_gpu,dig,6,22.594446
0.1,shared_gpu,face,6,256.022277
0.1,shared_gpu,ner,6,148.147381
0.1,dedicated_gpu,imc,6,22.916026
0.1,dedicated_gpu,dig,6,7.429501
0.1,dedicated_gpu,face,6,149.620071
0.1,dedicated_gpu,ner,6,48.434728
0.5,cpu,imc,6,2044.754324
0.5,cpu,dig,6,166.189636
0.5,cpu,face,6,5609.508364
0.5,cpu,ner,6,83.131868
0.5,shared_gpu,imc,6,20.652707
0.5,shared_gpu,dig,6,15.138819
0.5,shared_gpu,face,6,94.148688
0.5,shared_gpu,ner,6,44.719009
0.5,dedicated_gpu,imc,6,14.399452
0.5,dedicated_gpu,dig,6,7.115772
0.5,dedicated_gpu,face,6,96.865564
0.5,dedicated_gpu,ner,6,9.429311
1,cpu,imc,7,600.105172
1,cpu,dig,7,118.730254
1,cpu,face,7,1738.472781
1,cpu,ner,7,83.096812
1,shared_gpu,imc,7,11.50289
1,shared_gpu,dig,7,3.532977
1,shared_gpu,face,7,33.921883
1,shared_gpu,ner,7,23.325963
1,dedicated_gpu,imc,7,12.477551
1,dedicated_gpu,dig,7,5.646957
1,dedicated_gpu,face,7,37.863363
1,dedicated_gpu,ner,7,24.240751
0.25,cpu,imc,7,1689.88139
0.25,cpu,dig,7,195.786591
0.25,cpu,face,7,5183.490398
0.25,cpu,ner,7,159.209697
0.25,shared_gpu,imc,7,17.944943
0.25,shared_gpu,dig,7,10.043309
0.25,shared_gpu,face,7,97.73663
0.25,shared_gpu,ner,7,40.333423
0.25,dedicated_gpu,imc,7,23.351896
0.25,dedicated_gpu,dig,7,5.904611
0.25,dedicated_gpu,face,7,104.206378
0.25,dedicated_gpu,ner,7,7.390042
0.5,cpu,imc,7,1781.742212
0.5,cpu,dig,7,157.02621
0.5,cpu,face,7,5644.273889
0.5,cpu,ner,7,115.685267
0.5,shared_gpu,imc,7,17.720561
0.5,shared_gpu,dig,7,10.541658
0.5,shared_gpu,face,7,92.665932
0.5,shared_gpu,ner,7,44.036479
0.5,dedicated_gpu,imc,7,17.028875
0.5,dedicated_gpu,dig,7,3.431105
0.5,dedicated_gpu,face,7,74.550128
0.5,dedicated_gpu,ner,7,6.063055
0.1,cpu,imc,7,3356.174793
0.1,cpu,dig,7,358.293007
0.1,cpu,face,7,0
0.1,cpu,ner,7,140.960199
0.1,shared_gpu,imc,7,34.324623
0.1,shared_gpu,dig,7,18.9545
0.1,shared_gpu,face,7,185.759941
0.1,shared_gpu,ner,7,29.534543
0.1,dedicated_gpu,imc,7,31.554767
0.1,dedicated_gpu,dig,7,9.766318
0.1,dedicated_gpu,face,7,191.56923
0.1,dedicated_gpu,ner,7,52.748674
0.1,cpu,imc,8,3255.466596
0.1,cpu,dig,8,293.077306
0.1,cpu,face,8,0
0.1,cpu,ner,8,109.134092
0.1,shared_gpu,imc,8,35.553437
0.1,shared_gpu,dig,8,5.04283
0.1,shared_gpu,face,8,206.312515
0.1,shared_gpu,ner,8,24.753534
0.1,dedicated_gpu,imc,8,38.134492
0.1,dedicated_gpu,dig,8,4.401688
0.1,dedicated_gpu,face,8,145.422211
0.1,dedicated_gpu,ner,8,21.697567
1,cpu,imc,8,896.902226
1,cpu,dig,8,140.455769
1,cpu,face,8,2053.707358
1,cpu,ner,8,73.95756
1,shared_gpu,imc,8,13.032415
1,shared_gpu,dig,8,7.65672
1,shared_gpu,face,8,36.641806
1,shared_gpu,ner,8,14.512323
1,dedicated_gpu,imc,8,9.904043
1,dedicated_gpu,dig,8,6.719589
1,dedicated_gpu,face,8,40.043059
1,dedicated_gpu,ner,8,18.88697
0.25,cpu,imc,8,1607.960989
0.25,cpu,dig,8,152.563807
0.25,cpu,face,8,5076.646043
0.25,cpu,ner,8,97.452483
0.25,shared_gpu,imc,8,46.764197
0.25,shared_gpu,dig,8,19.424427
0.25,shared_gpu,face,8,110.301604
0.25,shared_gpu,ner,8,76.811297
0.25,dedicated_gpu,imc,8,25.07473
0.25,dedicated_gpu,dig,8,8.386667
0.25,dedicated_gpu,face,8,99.662723
0.25,dedicated_gpu,ner,8,3.909365
0.5,cpu,imc,8,1724.391297
0.5,cpu,dig,8,107.488765
0.5,cpu,face,8,5528.684248
0.5,cpu,ner,8,89.317459
0.5,shared_gpu,imc,8,15.324661
0.5,shared_gpu,dig,8,9.921452
0.5,shared_gpu,face,8,93.44809
0.5,shared_gpu,ner,8,41.340354
0.5,dedicated_gpu,imc,8,19.11275
0.5,dedicated_gpu,dig,8,9.581128
0.5,dedicated_gpu,face,8,0
0.5,dedicated_gpu,ner,8,0
0.1,cpu,imc,9,3194.988719
0.1,cpu,dig,9,289.350773
0.1,cpu,face,9,0
0.1,cpu,ner,9,70.560597
0.1,shared_gpu,imc,9,143.217261
0.1,shared_gpu,dig,9,27.438574
0.1,shared_gpu,face,9,240.957486
0.1,shared_gpu,ner,9,103.267568
0.1,dedicated_gpu,imc,9,30.342544
0.1,dedicated_gpu,dig,9,9.354402
0.1,dedicated_gpu,face,9,216.935008
0.1,dedicated_gpu,ner,9,212.202148
0.5,cpu,imc,9,1659.157889
0.5,cpu,dig,9,148.01475
0.5,cpu,face,9,5523.035945
0.5,cpu,ner,9,60.595038
0.5,shared_gpu,imc,9,29.041669
0.5,shared_gpu,dig,9,8.286074
0.5,shared_gpu,face,9,99.903847
0.5,shared_gpu,ner,9,49.52025
0.5,dedicated_gpu,imc,9,19.551769
0.5,dedicated_gpu,dig,9,5.969883
0.5,dedicated_gpu,face,9,97.07923
0.5,dedicated_gpu,ner,9,20.988234
1,cpu,imc,9,819.326243
1,cpu,dig,9,107.366636
1,cpu,face,9,2026.101148
1,cpu,ner,9,70.892
1,shared_gpu,imc,9,10.145899
1,shared_gpu,dig,9,8.23123
1,shared_gpu,face,9,33.281197
1,shared_gpu,ner,9,4.648711
1,dedicated_gpu,imc,9,15.397796
1,dedicated_gpu,dig,9,5.392608
1,dedicated_gpu,face,9,36.251779
1,dedicated_gpu,ner,9,8.242907
0.25,cpu,imc,9,1663.44643
0.25,cpu,dig,9,201.676494
0.25,cpu,face,9,5065.918558
0.25,cpu,ner,9,93.461442
0.25,shared_gpu,imc,9,19.307714
0.25,shared_gpu,dig,9,4.416767
0.25,shared_gpu,face,9,96.783553
0.25,shared_gpu,ner,9,73.652375
0.25,dedicated_gpu,imc,9,25.305667
0.25,dedicated_gpu,dig,9,8.564653
0.25,dedicated_gpu,face,9,89.354197
0.25,dedicated_gpu,ner,9,16.668341
1,cpu,imc,10,808.51427
1,cpu,dig,10,85.526389
1,cpu,face,10,2083.50043
1,cpu,ner,10,62.657145
1,shared_gpu,imc,10,18.412612
1,shared_gpu,dig,10,11.431406
1,shared_gpu,face,10,35.800345
1,shared_gpu,ner,10,10.001908
1,dedicated_gpu,imc,10,13.973715
1,dedicated_gpu,dig,10,7.123873
1,dedicated_gpu,face,10,36.81132
1,dedicated_gpu,ner,10,8.473017
0.1,cpu,imc,10,3449.908407
0.1,cpu,dig,10,316.743213
0.1,cpu,face,10,0
0.1,cpu,ner,10,83.115987
0.1,shared_gpu,imc,10,37.383678
0.1,shared_gpu,dig,10,7.226121
0.1,shared_gpu,face,10,193.447837
0.1,shared_gpu,ner,10,97.296398
0.1,dedicated_gpu,imc,10,51.919052
0.1,dedicated_gpu,dig,10,16.146258
0.1,dedicated_gpu,face,10,114.495981
0.1,dedicated_gpu,ner,10,13.924632
0.25,cpu,imc,10,1525.095261
0.25,cpu,dig,10,170.32719
0.25,cpu,face,10,5090.545444
0.25,cpu,ner,10,61.521739
0.25,shared_gpu,imc,10,26.025656
0.25,shared_gpu,dig,10,5.652431
0.25,shared_gpu,face,10,117.393674
0.25,shared_gpu,ner,10,28.445972
0.25,dedicated_gpu,imc,10,28.250785
0.25,dedicated_gpu,dig,10,9.505465
0.25,dedicated_gpu,face,10,102.896318
0.25,dedicated_gpu,ner,10,20.796574
0.5,cpu,imc,10,1932.280606
0.5,cpu,dig,10,152.501864
0.5,cpu,face,10,5740.430323
0.5,cpu,ner,10,86.785626
0.5,shared_gpu,imc,10,12.775512
0.5,shared_gpu,dig,10,3.316372
0.5,shared_gpu,face,10,91.934803
0.5,shared_gpu,ner,10,42.025754
0.5,dedicated_gpu,imc,10,28.962691
0.5,dedicated_gpu,dig,10,17.567869
0.5,dedicated_gpu,face,10,98.931294
0.5,dedicated_gpu,ner,10,24.8354
